*** SPICE deck for cell OneBitCam{sch} from library Project-1
*** Created on Sun Jul 02, 2023 09:43:46
*** Last revised on Sun Jul 02, 2023 10:49:45
*** Written on Sun Jul 02, 2023 10:49:49 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Project-1__SRAM FROM CELL SRAM{sch}
.SUBCKT Project-1__SRAM BL BLB Q QB RD vdd WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Q WL BL gnd nmos L=0.044U W=0.264U
Mnmos@1 BLB WL QB gnd nmos L=0.044U W=0.264U
Mnmos@2 net@28 Q BL gnd nmos L=0.044U W=0.132U
Mnmos@3 BLB QB net@28 gnd nmos L=0.044U W=0.132U
Mnmos@4 net@28 RD gnd gnd nmos L=0.044U W=0.198U
Mnmos@5 gnd QB Q gnd nmos L=0.044U W=0.066U
Mnmos@6 QB Q gnd gnd nmos L=0.044U W=0.066U
Mpmos@0 Q QB vdd vdd pmos L=0.044U W=0.066U
Mpmos@1 vdd Q QB vdd pmos L=0.044U W=0.066U
.ENDS Project-1__SRAM

.global gnd vdd

*** TOP LEVEL CELL: OneBitCam{sch}
Mnmos@0 Match net@19 net@15 gnd nmos L=0.044U W=0.044U
Mnmos@2 Match net@27 net@4 gnd nmos L=0.044U W=0.044U
Mnmos@3 net@4 CAM_Data gnd gnd nmos L=0.044U W=0.044U
Mnmos@4 net@15 net@4 gnd gnd nmos L=0.044U W=0.044U
Mpmos@0 net@15 net@27 Match vdd pmos L=0.044U W=0.044U
Mpmos@3 net@4 net@19 Match vdd pmos L=0.044U W=0.044U
Mpmos@4 vdd CAM_Data net@4 vdd pmos L=0.044U W=0.044U
Mpmos@5 vdd net@4 net@15 vdd pmos L=0.044U W=0.044U
XSRAM@1 BL BLB net@19 net@27 RD vdd WL Project-1__SRAM

* Spice Code nodes in cell cell 'OneBitCam{sch}'
vdd vdd 0 0.95
Vin_RL RL 0 PWL(0 0 10n 0 30n 0)
Vin_WL WL 0 PWL(0 0.95 20n 0.95 21n 0)
Vin_BL BL 0 PWL(0 0.95 20n 0.95 21n 0)
Vin_BLB BLB 0 PWL(0 0 20n 0 21n 0.95)
Vin_CAMDATA CAM_Data 0 PWL(0 0 20n 0 21n 0.95)
.tran 0 0.1us
.include C:\Program Files\LTC\LTspiceXVII\model\model.txt
.END
